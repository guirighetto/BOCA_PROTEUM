library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
 
entity <<ENTITY_NAME>> is
	port (<<IN_P>>: in <<type>>; <<OUT_P>>: out <<type>>);
end <<ENTITY_NAME>>;
 
architecture <<ARCH_TYPE>> of <<ENTITY_NAME>> is
  <<DECL_COMPONENTS>>
  <<DECL_SIGNALS>>
begin
  -- Commands.
  <<DECL_COMP_INSTANCES>>
end <<ARCH_TYPE>>;

