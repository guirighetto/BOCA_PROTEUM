-- Declaration of Components.\n
component <<COMPONENT_NAME>>\n
	port(<<ports_in>>: in <<type>>; <<ports_out>>: out <<type>>);\n
end component;\n
