-- Component instantiation and port mapping.\n
<<instance_name>>: <<COMPONENT_NAME>> port map(<<port1>>=><<portX>>, <<port2>>=><<portY>>);
